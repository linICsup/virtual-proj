`ifndef LIN_AHB_PKG_SV
`define LIN_AHB_PKG_SV

package lin_ahb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "lin_ahb_defines.svh"
  `include "lin_ahb_types.sv"
  `include "lin_ahb_configuration.sv"
  `include "lin_ahb_agent_configuration.sv"
  `include "lin_ahb_transaction.sv"
  `include "lin_ahb_sequencer.sv"
  `include "lin_ahb_driver.sv"
  `include "lin_ahb_monitor.sv"
  `include "lin_ahb_master_transaction.sv"
  `include "lin_ahb_master_driver.sv"
  `include "lin_ahb_master_monitor.sv"
  `include "lin_ahb_master_sequencer.sv"
  `include "lin_ahb_master_agent.sv"


  endpackage

`endif // LIN_AHB_PKG_SV
