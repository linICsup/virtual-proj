`ifndef LZC_AHBRAM_SEQ_LIB_SVH
`define LZC_AHBRAM_SEQ_LIB_SVH

`include "lzc_ahbram_base_virtual_sequencer.sv"
`include "lzc_ahbram_smoke_virt_seq.sv"

`endif
