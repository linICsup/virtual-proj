`ifndef LIN_AHB_IF_SV
`define LIN_AHB_IF_SV

interface lin_ahb_if;

endinterface

`endif // LIN_AHB_IF_SV
