`ifndef LZC_AHBRAM_TESTS_SVH
`define LZC_AHBRAM_TESTS_SVH

`include "lzc_ahbram_base_test.sv"
`include "lzc_ahbram_smoke_test.sv"

`endif // LZC_AHBRAM_TESTS_SVH
