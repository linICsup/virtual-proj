
module lzc_ahbram_tb;
import uvm_pkg::*;
`include "uvm_macros.svh"
import lzc_ahbram_pkg::*;

ahb_blockram_32 dut();

initial begin

end

endmodule
