`ifndef LIN_AHB_DEFINES_SVH
`define LIN_AHB_DEFINES_SVH

`define LIN_AHB_MAX_DATA_WIDTH 64
`define LIN_AHB_MAX_ADDR_WIDTH 32

`endif // LIN_AHB_DEFINES_SVH
