`ifndef LZC_AHBRAM_IF_SV
`define LZC_AHBRAM_IF_SV

interface lzc_ahbram_if;

endinterface


`endif // LZC_AHBRAM_IF_SV
