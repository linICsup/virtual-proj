`ifndef LZC_AHBRAM_PKG_SV
`define LZC_AHBRAM_PKG_SV

package lzc_ahbram_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
import lin_ahb_pkg::*;
endpackage
`endif  //LZC_AHBRAM_PKG_SV
